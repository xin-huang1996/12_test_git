module	test(
input	[3:0]	)